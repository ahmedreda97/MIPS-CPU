


library IEEE;
use IEEE.STD_LOGIC_1164.all;

package MyPackage is
component reg is

Generic(n:NATURAL :=4);
PORT(
I:IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
CLK,LD,INC,CLR :IN STD_LOGIC;
O:OUT STD_LOGIC_VECTOR(n-1 downto 0) );

end component;

component Decoder5x32 is

Port ( I : in  STD_LOGIC_VECTOR (4 downto 0);
           O : out  STD_LOGIC_VECTOR (31 downto 0));
end component;

component Mux2x1 is

Port (S : in  STD_LOGIC;
           I0 : in  STD_LOGIC;
           I1 : in  STD_LOGIC;
           O : out  STD_LOGIC);
end component;

component Mux4x1 is

 Port ( S : in  STD_LOGIC_VECTOR (1 downto 0);
           I0 : in  STD_LOGIC;
           I1 : in  STD_LOGIC;
           I2 : in  STD_LOGIC;
           I3 : in  STD_LOGIC;
           O : out  STD_LOGIC);

end component;

component Mux32x1 is

 Port ( S : in  STD_LOGIC_VECTOR (4 downto 0);
           I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,I16,I17,I18,I19,I20,I21,I22,I23,I24,I25,I26,I27,I28,I29,I30,I31 : in  STD_LOGIC_VECTOR (31 downto 0);
           O : out  STD_LOGIC_VECTOR (31 downto 0));

end component;

component OneBitALU is
Port (A : in  STD_LOGIC;
           B : in  STD_LOGIC;
			 SetLess:in std_logic;
			  AMuxop: in STD_LOGIC;
			  BMuxop : in STD_LOGIC;
			  MainMuxop : in STD_LOGIC_VECTOR(1 downto 0);
           CarryIn : in  STD_LOGIC;
           CarryOut : out  STD_LOGIC;
           Result : out  STD_LOGIC;
			  SetSum:out std_logic);
end component;
component Mux2x132bit is
 Port ( S : in  STD_LOGIC;
           I0 : in  STD_LOGIC_vector(31 downto 0);
           I1 : in  STD_LOGIC_vector(31 downto 0);
           O : out  STD_LOGIC_vector(31 downto 0));
end component;

end MyPackage;

package body MyPackage is


 
end MyPackage;
